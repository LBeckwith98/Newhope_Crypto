`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Virginia Tech
// Engineer: Luke Beckwith
// 
// Create Date: 05/07/2019 10:37:11 PM
// Module Name: omega
// Project Name:  NTT
// Description: Given the bf_num and layer, this determines what
//  omega should be the input to the butterfly module
//////////////////////////////////////////////////////////////////////////////////


module omega_lut(
    input clk,
    input [3:0] layer_num,
    input [7:0] bf_num,
    input inverse,
    output reg [15:0] omega_out
    );

    wire [7:0] omega_sel;
    assign omega_sel = (layer_num == 0) ? bf_num & 8'hFF :
                        (layer_num == 1) ? bf_num & 8'h7F :
                        (layer_num == 2) ? bf_num & 8'h3F :
                        (layer_num == 3) ? bf_num & 8'h1F :
                        (layer_num == 4) ? bf_num & 8'h0F :
                        (layer_num == 5) ? bf_num & 8'h07 :
                        (layer_num == 6) ? bf_num & 8'h03 :
                        (layer_num == 7) ? bf_num & 8'h01 : 8'h00;

    always @(posedge clk) begin
        if (inverse == 0) begin
            case (omega_sel)
               8'd0: omega_out = 16'd4075;
               8'd1: omega_out = 16'd5315;
               8'd2: omega_out = 16'd7965;
               8'd3: omega_out = 16'd7373;
               8'd4: omega_out = 16'd522;
               8'd5: omega_out = 16'd10120;
               8'd6: omega_out = 16'd9027;
               8'd7: omega_out = 16'd5079;
               8'd8: omega_out = 16'd2344;
               8'd9: omega_out = 16'd1278;
               8'd10: omega_out = 16'd1973;
               8'd11: omega_out = 16'd5574;
               8'd12: omega_out = 16'd1018;
               8'd13: omega_out = 16'd6364;
               8'd14: omega_out = 16'd11248;
               8'd15: omega_out = 16'd8775;
               8'd16: omega_out = 16'd7500;
               8'd17: omega_out = 16'd7822;
               8'd18: omega_out = 16'd5537;
               8'd19: omega_out = 16'd4749;
               8'd20: omega_out = 16'd8500;
               8'd21: omega_out = 16'd12142;
               8'd22: omega_out = 16'd5456;
               8'd23: omega_out = 16'd7840;
               8'd24: omega_out = 16'd5445;
               8'd25: omega_out = 16'd3860;
               8'd26: omega_out = 16'd4536;
               8'd27: omega_out = 16'd11239;
               8'd28: omega_out = 16'd6171;
               8'd29: omega_out = 16'd8471;
               8'd30: omega_out = 16'd2683;
               8'd31: omega_out = 16'd11099;
               8'd32: omega_out = 16'd10561;
               8'd33: omega_out = 16'd400;
               8'd34: omega_out = 16'd6137;
               8'd35: omega_out = 16'd7341;
               8'd36: omega_out = 16'd5415;
               8'd37: omega_out = 16'd8646;
               8'd38: omega_out = 16'd6136;
               8'd39: omega_out = 16'd5862;
               8'd40: omega_out = 16'd5529;
               8'd41: omega_out = 16'd5206;
               8'd42: omega_out = 16'd56;
               8'd43: omega_out = 16'd9090;
               8'd44: omega_out = 16'd8724;
               8'd45: omega_out = 16'd11635;
               8'd46: omega_out = 16'd1702;
               8'd47: omega_out = 16'd10302;
               8'd48: omega_out = 16'd5339;
               8'd49: omega_out = 16'd6843;
               8'd50: omega_out = 16'd6093;
               8'd51: omega_out = 16'd3710;
               8'd52: omega_out = 16'd316;
               8'd53: omega_out = 16'd382;
               8'd54: omega_out = 16'd11821;
               8'd55: omega_out = 16'd8301;
               8'd56: omega_out = 16'd10930;
               8'd57: omega_out = 16'd5435;
               8'd58: omega_out = 16'd11035;
               8'd59: omega_out = 16'd973;
               8'd60: omega_out = 16'd8291;
               8'd61: omega_out = 16'd10256;
               8'd62: omega_out = 16'd8410;
               8'd63: omega_out = 16'd1922;
               8'd64: omega_out = 16'd12097;
               8'd65: omega_out = 16'd10968;
               8'd66: omega_out = 16'd10240;
               8'd67: omega_out = 16'd4912;
               8'd68: omega_out = 16'd4698;
               8'd69: omega_out = 16'd5057;
               8'd70: omega_out = 16'd7509;
               8'd71: omega_out = 16'd8844;
               8'd72: omega_out = 16'd8807;
               8'd73: omega_out = 16'd11502;
               8'd74: omega_out = 16'd5468;
               8'd75: omega_out = 16'd1010;
               8'd76: omega_out = 16'd9162;
               8'd77: omega_out = 16'd8120;
               8'd78: omega_out = 16'd2920;
               8'd79: omega_out = 16'd5241;
               8'd80: omega_out = 16'd6055;
               8'd81: omega_out = 16'd8953;
               8'd82: omega_out = 16'd677;
               8'd83: omega_out = 16'd5874;
               8'd84: omega_out = 16'd2766;
               8'd85: omega_out = 16'd10966;
               8'd86: omega_out = 16'd12237;
               8'd87: omega_out = 16'd9115;
               8'd88: omega_out = 16'd12138;
               8'd89: omega_out = 16'd10162;
               8'd90: omega_out = 16'd3957;
               8'd91: omega_out = 16'd2839;
               8'd92: omega_out = 16'd6383;
               8'd93: omega_out = 16'd2505;
               8'd94: omega_out = 16'd11858;
               8'd95: omega_out = 16'd1579;
               8'd96: omega_out = 16'd9026;
               8'd97: omega_out = 16'd3600;
               8'd98: omega_out = 16'd6077;
               8'd99: omega_out = 16'd4624;
               8'd100: omega_out = 16'd11868;
               8'd101: omega_out = 16'd4080;
               8'd102: omega_out = 16'd6068;
               8'd103: omega_out = 16'd3602;
               8'd104: omega_out = 16'd605;
               8'd105: omega_out = 16'd9987;
               8'd106: omega_out = 16'd504;
               8'd107: omega_out = 16'd8076;
               8'd108: omega_out = 16'd4782;
               8'd109: omega_out = 16'd6403;
               8'd110: omega_out = 16'd3029;
               8'd111: omega_out = 16'd6695;
               8'd112: omega_out = 16'd11184;
               8'd113: omega_out = 16'd142;
               8'd114: omega_out = 16'd5681;
               8'd115: omega_out = 16'd8812;
               8'd116: omega_out = 16'd2844;
               8'd117: omega_out = 16'd3438;
               8'd118: omega_out = 16'd8077;
               8'd119: omega_out = 16'd975;
               8'd120: omega_out = 16'd58;
               8'd121: omega_out = 16'd12048;
               8'd122: omega_out = 16'd1003;
               8'd123: omega_out = 16'd8757;
               8'd124: omega_out = 16'd885;
               8'd125: omega_out = 16'd6281;
               8'd126: omega_out = 16'd1956;
               8'd127: omega_out = 16'd5009;
               8'd128: omega_out = 16'd12225;
               8'd129: omega_out = 16'd3656;
               8'd130: omega_out = 16'd11606;
               8'd131: omega_out = 16'd9830;
               8'd132: omega_out = 16'd1566;
               8'd133: omega_out = 16'd5782;
               8'd134: omega_out = 16'd2503;
               8'd135: omega_out = 16'd2948;
               8'd136: omega_out = 16'd7032;
               8'd137: omega_out = 16'd3834;
               8'd138: omega_out = 16'd5919;
               8'd139: omega_out = 16'd4433;
               8'd140: omega_out = 16'd3054;
               8'd141: omega_out = 16'd6803;
               8'd142: omega_out = 16'd9166;
               8'd143: omega_out = 16'd1747;
               8'd144: omega_out = 16'd10211;
               8'd145: omega_out = 16'd11177;
               8'd146: omega_out = 16'd4322;
               8'd147: omega_out = 16'd1958;
               8'd148: omega_out = 16'd922;
               8'd149: omega_out = 16'd11848;
               8'd150: omega_out = 16'd4079;
               8'd151: omega_out = 16'd11231;
               8'd152: omega_out = 16'd4046;
               8'd153: omega_out = 16'd11580;
               8'd154: omega_out = 16'd1319;
               8'd155: omega_out = 16'd9139;
               8'd156: omega_out = 16'd6224;
               8'd157: omega_out = 16'd835;
               8'd158: omega_out = 16'd8049;
               8'd159: omega_out = 16'd8719;
               8'd160: omega_out = 16'd7105;
               8'd161: omega_out = 16'd1200;
               8'd162: omega_out = 16'd6122;
               8'd163: omega_out = 16'd9734;
               8'd164: omega_out = 16'd3956;
               8'd165: omega_out = 16'd1360;
               8'd166: omega_out = 16'd6119;
               8'd167: omega_out = 16'd5297;
               8'd168: omega_out = 16'd4298;
               8'd169: omega_out = 16'd3329;
               8'd170: omega_out = 16'd168;
               8'd171: omega_out = 16'd2692;
               8'd172: omega_out = 16'd1594;
               8'd173: omega_out = 16'd10327;
               8'd174: omega_out = 16'd5106;
               8'd175: omega_out = 16'd6328;
               8'd176: omega_out = 16'd3728;
               8'd177: omega_out = 16'd8240;
               8'd178: omega_out = 16'd5990;
               8'd179: omega_out = 16'd11130;
               8'd180: omega_out = 16'd948;
               8'd181: omega_out = 16'd1146;
               8'd182: omega_out = 16'd10885;
               8'd183: omega_out = 16'd325;
               8'd184: omega_out = 16'd8212;
               8'd185: omega_out = 16'd4016;
               8'd186: omega_out = 16'd8527;
               8'd187: omega_out = 16'd2919;
               8'd188: omega_out = 16'd295;
               8'd189: omega_out = 16'd6190;
               8'd190: omega_out = 16'd652;
               8'd191: omega_out = 16'd5766;
               8'd192: omega_out = 16'd11713;
               8'd193: omega_out = 16'd8326;
               8'd194: omega_out = 16'd6142;
               8'd195: omega_out = 16'd2447;
               8'd196: omega_out = 16'd1805;
               8'd197: omega_out = 16'd2882;
               8'd198: omega_out = 16'd10238;
               8'd199: omega_out = 16'd1954;
               8'd200: omega_out = 16'd1843;
               8'd201: omega_out = 16'd9928;
               8'd202: omega_out = 16'd4115;
               8'd203: omega_out = 16'd3030;
               8'd204: omega_out = 16'd2908;
               8'd205: omega_out = 16'd12071;
               8'd206: omega_out = 16'd8760;
               8'd207: omega_out = 16'd3434;
               8'd208: omega_out = 16'd5876;
               8'd209: omega_out = 16'd2281;
               8'd210: omega_out = 16'd2031;
               8'd211: omega_out = 16'd5333;
               8'd212: omega_out = 16'd8298;
               8'd213: omega_out = 16'd8320;
               8'd214: omega_out = 16'd12133;
               8'd215: omega_out = 16'd2767;
               8'd216: omega_out = 16'd11836;
               8'd217: omega_out = 16'd5908;
               8'd218: omega_out = 16'd11871;
               8'd219: omega_out = 16'd8517;
               8'd220: omega_out = 16'd6860;
               8'd221: omega_out = 16'd7515;
               8'd222: omega_out = 16'd10996;
               8'd223: omega_out = 16'd4737;
               8'd224: omega_out = 16'd2500;
               8'd225: omega_out = 16'd10800;
               8'd226: omega_out = 16'd5942;
               8'd227: omega_out = 16'd1583;
               8'd228: omega_out = 16'd11026;
               8'd229: omega_out = 16'd12240;
               8'd230: omega_out = 16'd5915;
               8'd231: omega_out = 16'd10806;
               8'd232: omega_out = 16'd1815;
               8'd233: omega_out = 16'd5383;
               8'd234: omega_out = 16'd1512;
               8'd235: omega_out = 16'd11939;
               8'd236: omega_out = 16'd2057;
               8'd237: omega_out = 16'd6920;
               8'd238: omega_out = 16'd9087;
               8'd239: omega_out = 16'd7796;
               8'd240: omega_out = 16'd8974;
               8'd241: omega_out = 16'd426;
               8'd242: omega_out = 16'd4754;
               8'd243: omega_out = 16'd1858;
               8'd244: omega_out = 16'd8532;
               8'd245: omega_out = 16'd10314;
               8'd246: omega_out = 16'd11942;
               8'd247: omega_out = 16'd2925;
               8'd248: omega_out = 16'd174;
               8'd249: omega_out = 16'd11566;
               8'd250: omega_out = 16'd3009;
               8'd251: omega_out = 16'd1693;
               8'd252: omega_out = 16'd2655;
               8'd253: omega_out = 16'd6554;
               8'd254: omega_out = 16'd5868;
               8'd255: omega_out = 16'd2738;
            endcase
            end
        else begin
            case (omega_sel)
               8'd0: omega_out = 16'd4075;
               8'd1: omega_out = 16'd6974;
               8'd2: omega_out = 16'd4916;
               8'd3: omega_out = 16'd4324;
               8'd4: omega_out = 16'd7210;
               8'd5: omega_out = 16'd3262;
               8'd6: omega_out = 16'd2169;
               8'd7: omega_out = 16'd11767;
               8'd8: omega_out = 16'd3514;
               8'd9: omega_out = 16'd1041;
               8'd10: omega_out = 16'd5925;
               8'd11: omega_out = 16'd11271;
               8'd12: omega_out = 16'd6715;
               8'd13: omega_out = 16'd10316;
               8'd14: omega_out = 16'd11011;
               8'd15: omega_out = 16'd9945;
               8'd16: omega_out = 16'd1190;
               8'd17: omega_out = 16'd9606;
               8'd18: omega_out = 16'd3818;
               8'd19: omega_out = 16'd6118;
               8'd20: omega_out = 16'd1050;
               8'd21: omega_out = 16'd7753;
               8'd22: omega_out = 16'd8429;
               8'd23: omega_out = 16'd6844;
               8'd24: omega_out = 16'd4449;
               8'd25: omega_out = 16'd6833;
               8'd26: omega_out = 16'd147;
               8'd27: omega_out = 16'd3789;
               8'd28: omega_out = 16'd7540;
               8'd29: omega_out = 16'd6752;
               8'd30: omega_out = 16'd4467;
               8'd31: omega_out = 16'd4789;
               8'd32: omega_out = 16'd10367;
               8'd33: omega_out = 16'd3879;
               8'd34: omega_out = 16'd2033;
               8'd35: omega_out = 16'd3998;
               8'd36: omega_out = 16'd11316;
               8'd37: omega_out = 16'd1254;
               8'd38: omega_out = 16'd6854;
               8'd39: omega_out = 16'd1359;
               8'd40: omega_out = 16'd3988;
               8'd41: omega_out = 16'd468;
               8'd42: omega_out = 16'd11907;
               8'd43: omega_out = 16'd11973;
               8'd44: omega_out = 16'd8579;
               8'd45: omega_out = 16'd6196;
               8'd46: omega_out = 16'd5446;
               8'd47: omega_out = 16'd6950;
               8'd48: omega_out = 16'd1987;
               8'd49: omega_out = 16'd10587;
               8'd50: omega_out = 16'd654;
               8'd51: omega_out = 16'd3565;
               8'd52: omega_out = 16'd3199;
               8'd53: omega_out = 16'd12233;
               8'd54: omega_out = 16'd7083;
               8'd55: omega_out = 16'd6760;
               8'd56: omega_out = 16'd6427;
               8'd57: omega_out = 16'd6153;
               8'd58: omega_out = 16'd3643;
               8'd59: omega_out = 16'd6874;
               8'd60: omega_out = 16'd4948;
               8'd61: omega_out = 16'd6152;
               8'd62: omega_out = 16'd11889;
               8'd63: omega_out = 16'd1728;
               8'd64: omega_out = 16'd7280;
               8'd65: omega_out = 16'd10333;
               8'd66: omega_out = 16'd6008;
               8'd67: omega_out = 16'd11404;
               8'd68: omega_out = 16'd3532;
               8'd69: omega_out = 16'd11286;
               8'd70: omega_out = 16'd241;
               8'd71: omega_out = 16'd12231;
               8'd72: omega_out = 16'd11314;
               8'd73: omega_out = 16'd4212;
               8'd74: omega_out = 16'd8851;
               8'd75: omega_out = 16'd9445;
               8'd76: omega_out = 16'd3477;
               8'd77: omega_out = 16'd6608;
               8'd78: omega_out = 16'd12147;
               8'd79: omega_out = 16'd1105;
               8'd80: omega_out = 16'd5594;
               8'd81: omega_out = 16'd9260;
               8'd82: omega_out = 16'd5886;
               8'd83: omega_out = 16'd7507;
               8'd84: omega_out = 16'd4213;
               8'd85: omega_out = 16'd11785;
               8'd86: omega_out = 16'd2302;
               8'd87: omega_out = 16'd11684;
               8'd88: omega_out = 16'd8687;
               8'd89: omega_out = 16'd6221;
               8'd90: omega_out = 16'd8209;
               8'd91: omega_out = 16'd421;
               8'd92: omega_out = 16'd7665;
               8'd93: omega_out = 16'd6212;
               8'd94: omega_out = 16'd8689;
               8'd95: omega_out = 16'd3263;
               8'd96: omega_out = 16'd10710;
               8'd97: omega_out = 16'd431;
               8'd98: omega_out = 16'd9784;
               8'd99: omega_out = 16'd5906;
               8'd100: omega_out = 16'd9450;
               8'd101: omega_out = 16'd8332;
               8'd102: omega_out = 16'd2127;
               8'd103: omega_out = 16'd151;
               8'd104: omega_out = 16'd3174;
               8'd105: omega_out = 16'd52;
               8'd106: omega_out = 16'd1323;
               8'd107: omega_out = 16'd9523;
               8'd108: omega_out = 16'd6415;
               8'd109: omega_out = 16'd11612;
               8'd110: omega_out = 16'd3336;
               8'd111: omega_out = 16'd6234;
               8'd112: omega_out = 16'd7048;
               8'd113: omega_out = 16'd9369;
               8'd114: omega_out = 16'd4169;
               8'd115: omega_out = 16'd3127;
               8'd116: omega_out = 16'd11279;
               8'd117: omega_out = 16'd6821;
               8'd118: omega_out = 16'd787;
               8'd119: omega_out = 16'd3482;
               8'd120: omega_out = 16'd3445;
               8'd121: omega_out = 16'd4780;
               8'd122: omega_out = 16'd7232;
               8'd123: omega_out = 16'd7591;
               8'd124: omega_out = 16'd7377;
               8'd125: omega_out = 16'd2049;
               8'd126: omega_out = 16'd1321;
               8'd127: omega_out = 16'd192;
               8'd128: omega_out = 16'd9551;
               8'd129: omega_out = 16'd6421;
               8'd130: omega_out = 16'd5735;
               8'd131: omega_out = 16'd9634;
               8'd132: omega_out = 16'd10596;
               8'd133: omega_out = 16'd9280;
               8'd134: omega_out = 16'd723;
               8'd135: omega_out = 16'd12115;
               8'd136: omega_out = 16'd9364;
               8'd137: omega_out = 16'd347;
               8'd138: omega_out = 16'd1975;
               8'd139: omega_out = 16'd3757;
               8'd140: omega_out = 16'd10431;
               8'd141: omega_out = 16'd7535;
               8'd142: omega_out = 16'd11863;
               8'd143: omega_out = 16'd3315;
               8'd144: omega_out = 16'd4493;
               8'd145: omega_out = 16'd3202;
               8'd146: omega_out = 16'd5369;
               8'd147: omega_out = 16'd10232;
               8'd148: omega_out = 16'd350;
               8'd149: omega_out = 16'd10777;
               8'd150: omega_out = 16'd6906;
               8'd151: omega_out = 16'd10474;
               8'd152: omega_out = 16'd1483;
               8'd153: omega_out = 16'd6374;
               8'd154: omega_out = 16'd49;
               8'd155: omega_out = 16'd1263;
               8'd156: omega_out = 16'd10706;
               8'd157: omega_out = 16'd6347;
               8'd158: omega_out = 16'd1489;
               8'd159: omega_out = 16'd9789;
               8'd160: omega_out = 16'd7552;
               8'd161: omega_out = 16'd1293;
               8'd162: omega_out = 16'd4774;
               8'd163: omega_out = 16'd5429;
               8'd164: omega_out = 16'd3772;
               8'd165: omega_out = 16'd418;
               8'd166: omega_out = 16'd6381;
               8'd167: omega_out = 16'd453;
               8'd168: omega_out = 16'd9522;
               8'd169: omega_out = 16'd156;
               8'd170: omega_out = 16'd3969;
               8'd171: omega_out = 16'd3991;
               8'd172: omega_out = 16'd6956;
               8'd173: omega_out = 16'd10258;
               8'd174: omega_out = 16'd10008;
               8'd175: omega_out = 16'd6413;
               8'd176: omega_out = 16'd8855;
               8'd177: omega_out = 16'd3529;
               8'd178: omega_out = 16'd218;
               8'd179: omega_out = 16'd9381;
               8'd180: omega_out = 16'd9259;
               8'd181: omega_out = 16'd8174;
               8'd182: omega_out = 16'd2361;
               8'd183: omega_out = 16'd10446;
               8'd184: omega_out = 16'd10335;
               8'd185: omega_out = 16'd2051;
               8'd186: omega_out = 16'd9407;
               8'd187: omega_out = 16'd10484;
               8'd188: omega_out = 16'd9842;
               8'd189: omega_out = 16'd6147;
               8'd190: omega_out = 16'd3963;
               8'd191: omega_out = 16'd576;
               8'd192: omega_out = 16'd6523;
               8'd193: omega_out = 16'd11637;
               8'd194: omega_out = 16'd6099;
               8'd195: omega_out = 16'd11994;
               8'd196: omega_out = 16'd9370;
               8'd197: omega_out = 16'd3762;
               8'd198: omega_out = 16'd8273;
               8'd199: omega_out = 16'd4077;
               8'd200: omega_out = 16'd11964;
               8'd201: omega_out = 16'd1404;
               8'd202: omega_out = 16'd11143;
               8'd203: omega_out = 16'd11341;
               8'd204: omega_out = 16'd1159;
               8'd205: omega_out = 16'd6299;
               8'd206: omega_out = 16'd4049;
               8'd207: omega_out = 16'd8561;
               8'd208: omega_out = 16'd5961;
               8'd209: omega_out = 16'd7183;
               8'd210: omega_out = 16'd1962;
               8'd211: omega_out = 16'd10695;
               8'd212: omega_out = 16'd9597;
               8'd213: omega_out = 16'd12121;
               8'd214: omega_out = 16'd8960;
               8'd215: omega_out = 16'd7991;
               8'd216: omega_out = 16'd6992;
               8'd217: omega_out = 16'd6170;
               8'd218: omega_out = 16'd10929;
               8'd219: omega_out = 16'd8333;
               8'd220: omega_out = 16'd2555;
               8'd221: omega_out = 16'd6167;
               8'd222: omega_out = 16'd11089;
               8'd223: omega_out = 16'd5184;
               8'd224: omega_out = 16'd3570;
               8'd225: omega_out = 16'd4240;
               8'd226: omega_out = 16'd11454;
               8'd227: omega_out = 16'd6065;
               8'd228: omega_out = 16'd3150;
               8'd229: omega_out = 16'd10970;
               8'd230: omega_out = 16'd709;
               8'd231: omega_out = 16'd8243;
               8'd232: omega_out = 16'd1058;
               8'd233: omega_out = 16'd8210;
               8'd234: omega_out = 16'd441;
               8'd235: omega_out = 16'd11367;
               8'd236: omega_out = 16'd10331;
               8'd237: omega_out = 16'd7967;
               8'd238: omega_out = 16'd1112;
               8'd239: omega_out = 16'd2078;
               8'd240: omega_out = 16'd10542;
               8'd241: omega_out = 16'd3123;
               8'd242: omega_out = 16'd5486;
               8'd243: omega_out = 16'd9235;
               8'd244: omega_out = 16'd7856;
               8'd245: omega_out = 16'd6370;
               8'd246: omega_out = 16'd8455;
               8'd247: omega_out = 16'd5257;
               8'd248: omega_out = 16'd9341;
               8'd249: omega_out = 16'd9786;
               8'd250: omega_out = 16'd6507;
               8'd251: omega_out = 16'd10723;
               8'd252: omega_out = 16'd2459;
               8'd253: omega_out = 16'd683;
               8'd254: omega_out = 16'd8633;
               8'd255: omega_out = 16'd64;
            endcase
        end   
    end
       
endmodule
