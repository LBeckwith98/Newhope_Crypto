`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Create Date: 05/08/2019 03:18:03 PM
// Module Name: poly_ram
// Project Name:  NTT
// Description: Vivado BRAM block. 
// (https://www.xilinx.com/support/documentation/sw_manuals/xilinx2018_3/ug901-vivado-synthesis.pdf)
// Page 122
//////////////////////////////////////////////////////////////////////////////////


module poly_ram (clka,clkb,ena,enb,wea,web,addra,addrb,dia,dib,doa,dob);
    parameter FILENAME = "";

    input clka, clkb, ena, enb, wea, web;
    input [10:0] addra, addrb;
    input [15:0] dia, dib;
    output [15:0] doa, dob;
    reg [15:0] ram [2047:0];
    reg [15:0] doa, dob;
        
    // addr a logic
    always @(posedge clka)
    begin
        if (ena)
        begin
            if (wea)
                ram[addra] <= dia;
            doa <= ram[addra];
        end
    end
    
    // addrb logic
    always @(posedge clkb)
        begin
        if (enb)
        begin
            if (web)
                ram[addrb] <= dib;
            dob <= ram[addrb];
        end
    end
    
    // initialize top of RAM with gammas_inv_montgomery
    initial begin
      if (FILENAME != "") begin
        $readmemh(FILENAME, ram);
      end
    end
       /*if (INVERSE_GAMMAS == 1'b1) begin
        ram[0] = 16'h0200;
        ram[1] = 16'h0F68;
        ram[2] = 16'h10AB;
        ram[3] = 16'h1523;
        ram[4] = 16'h258F;
        ram[5] = 16'h170C;
        ram[6] = 16'h0C85;
        ram[7] = 16'h17AF;
        ram[8] = 16'h242D;
        ram[9] = 16'h07E5;
        ram[10] = 16'h0C0F;
        ram[11] = 16'h12A2;
        ram[12] = 16'h0405;
        ram[13] = 16'h0636;
        ram[14] = 16'h0157;
        ram[15] = 16'h0212;
        ram[16] = 16'h2073;
        ram[17] = 16'h10B1;
        ram[18] = 16'h0AD1;
        ram[19] = 16'h2591;
        ram[20] = 16'h039B;
        ram[21] = 16'h1C86;
        ram[22] = 16'h1134;
        ram[23] = 16'h0982;
        ram[24] = 16'h05BC;
        ram[25] = 16'h232C;
        ram[26] = 16'h21EA;
        ram[27] = 16'h2BBA;
        ram[28] = 16'h0B4E;
        ram[29] = 16'h2E94;
        ram[30] = 16'h13C5;
        ram[31] = 16'h1F87;
        ram[32] = 16'h0697;
        ram[33] = 16'h2A83;
        ram[34] = 16'h2233;
        ram[35] = 16'h1E2C;
        ram[36] = 16'h2B67;
        ram[37] = 16'h1A0F;
        ram[38] = 16'h1E78;
        ram[39] = 16'h18B0;
        ram[40] = 16'h0A28;
        ram[41] = 16'h183B;
        ram[42] = 16'h1363;
        ram[43] = 16'h1814;
        ram[44] = 16'h2677;
        ram[45] = 16'h1807;
        ram[46] = 16'h2CD3;
        ram[47] = 16'h2803;
        ram[48] = 16'h0EF1;
        ram[49] = 16'h2D57;
        ram[50] = 16'h04FB;
        ram[51] = 16'h0F1D;
        ram[52] = 16'h01A9;
        ram[53] = 16'h150A;
        ram[54] = 16'h108E;
        ram[55] = 16'h2704;
        ram[56] = 16'h1585;
        ram[57] = 16'h2D02;
        ram[58] = 16'h272D;
        ram[59] = 16'h1F01;
        ram[60] = 16'h0D0F;
        ram[61] = 16'h1A56;
        ram[62] = 16'h245B;
        ram[63] = 16'h28C8;
        ram[64] = 16'h2C1F;
        ram[65] = 16'h0D98;
        ram[66] = 16'h0EB5;
        ram[67] = 16'h0488;
        ram[68] = 16'h04E7;
        ram[69] = 16'h1183;
        ram[70] = 16'h21A3;
        ram[71] = 16'h25D7;
        ram[72] = 16'h2B37;
        ram[73] = 16'h0C9D;
        ram[74] = 16'h1E68;
        ram[75] = 16'h2435;
        ram[76] = 16'h1A23;
        ram[77] = 16'h1C12;
        ram[78] = 16'h28B7;
        ram[79] = 16'h295C;
        ram[80] = 16'h2D93;
        ram[81] = 16'h2DCA;
        ram[82] = 16'h0F31;
        ram[83] = 16'h2F44;
        ram[84] = 16'h2511;
        ram[85] = 16'h2FC2;
        ram[86] = 16'h0C5B;
        ram[87] = 16'h2FEC;
        ram[88] = 16'h241F;
        ram[89] = 16'h2FFA;
        ram[90] = 16'h2C0B;
        ram[91] = 16'h0FFE;
        ram[92] = 16'h2EAF;
        ram[93] = 16'h1555;
        ram[94] = 16'h1F90;
        ram[95] = 16'h271D;
        ram[96] = 16'h2A86;
        ram[97] = 16'h1D0A;
        ram[98] = 16'h1E2D;
        ram[99] = 16'h09AE;
        ram[100] = 16'h0A0F;
        ram[101] = 16'h033A;
        ram[102] = 16'h235B;
        ram[103] = 16'h2114;
        ram[104] = 16'h0BC9;
        ram[105] = 16'h1B07;
        ram[106] = 16'h13EE;
        ram[107] = 16'h2903;
        ram[108] = 16'h16A5;
        ram[109] = 16'h1DAC;
        ram[110] = 16'h278D;
        ram[111] = 16'h09E4;
        ram[112] = 16'h0D2F;
        ram[113] = 16'h034C;
        ram[114] = 16'h0465;
        ram[115] = 16'h211A;
        ram[116] = 16'h0177;
        ram[117] = 16'h1B09;
        ram[118] = 16'h007D;
        ram[119] = 16'h0903;
        ram[120] = 16'h102A;
        ram[121] = 16'h0301;
        ram[122] = 16'h2564;
        ram[123] = 16'h2101;
        ram[124] = 16'h1C77;
        ram[125] = 16'h2B01;
        ram[126] = 16'h097D;
        ram[127] = 16'h1E56;
        ram[128] = 16'h132A;
        ram[129] = 16'h1A1D;
        ram[130] = 16'h2664;
        ram[131] = 16'h28B5;
        ram[132] = 16'h0CCC;
        ram[133] = 16'h1D92;
        ram[134] = 16'h0444;
        ram[135] = 16'h29DC;
        ram[136] = 16'h016C;
        ram[137] = 16'h0DF4;
        ram[138] = 16'h207A;
        ram[139] = 16'h14A7;
        ram[140] = 16'h2AD4;
        ram[141] = 16'h26E3;
        ram[142] = 16'h1E47;
        ram[143] = 16'h2CF7;
        ram[144] = 16'h1A18;
        ram[145] = 16'h0EFD;
        ram[146] = 16'h18B3;
        ram[147] = 16'h04FF;
        ram[148] = 16'h183C;
        ram[149] = 16'h21AB;
        ram[150] = 16'h0814;
        ram[151] = 16'h0B39;
        ram[152] = 16'h22B2;
        ram[153] = 16'h13BE;
        ram[154] = 16'h1B91;
        ram[155] = 16'h1695;
        ram[156] = 16'h2931;
        ram[157] = 16'h0787;
        ram[158] = 16'h0DBB;
        ram[159] = 16'h2283;
        ram[160] = 16'h1494;
        ram[161] = 16'h0B81;
        ram[162] = 16'h06DC;
        ram[163] = 16'h13D6;
        ram[164] = 16'h224A;
        ram[165] = 16'h169D;
        ram[166] = 16'h0B6E;
        ram[167] = 16'h178A;
        ram[168] = 16'h23D0;
        ram[169] = 16'h17D9;
        ram[170] = 16'h0BF0;
        ram[171] = 16'h07F3;
        ram[172] = 16'h13FB;
        ram[173] = 16'h22A7;
        ram[174] = 16'h06A9;
        ram[175] = 16'h0B8D;
        ram[176] = 16'h2239;
        ram[177] = 16'h13DA;
        ram[178] = 16'h2B69;
        ram[179] = 16'h069E;
        ram[180] = 16'h2E79;
        ram[181] = 16'h1235;
        ram[182] = 16'h1F7E;
        ram[183] = 16'h1612;
        ram[184] = 16'h2A80;
        ram[185] = 16'h275C;
        ram[186] = 16'h1E2B;
        ram[187] = 16'h1D1F;
        ram[188] = 16'h2A0F;
        ram[189] = 16'h09B5;
        ram[190] = 16'h0E05;
        ram[191] = 16'h233D;
        ram[192] = 16'h24AD;
        ram[193] = 16'h0BBF;
        ram[194] = 16'h1C3A;
        ram[195] = 16'h23EB;
        ram[196] = 16'h1969;
        ram[197] = 16'h0BF9;
        ram[198] = 16'h2879;
        ram[199] = 16'h13FE;
        ram[200] = 16'h1D7E;
        ram[201] = 16'h06AA;
        ram[202] = 16'h19D5;
        ram[203] = 16'h1239;
        ram[204] = 16'h289D;
        ram[205] = 16'h0613;
        ram[206] = 16'h1D8A;
        ram[207] = 16'h2207;
        ram[208] = 16'h19D9;
        ram[209] = 16'h1B58;
        ram[210] = 16'h189E;
        ram[211] = 16'h291E;
        ram[212] = 16'h1835;
        ram[213] = 16'h1DB5;
        ram[214] = 16'h1812;
        ram[215] = 16'h09E7;
        ram[216] = 16'h0806;
        ram[217] = 16'h034D;
        ram[218] = 16'h12AD;
        ram[219] = 16'h111A;
        ram[220] = 16'h163A;
        ram[221] = 16'h25B4;
        ram[222] = 16'h1769;
        ram[223] = 16'h2C92;
        ram[224] = 16'h17CE;
        ram[225] = 16'h2EDC;
        ram[226] = 16'h27F0;
        ram[227] = 16'h1F9F;
        ram[228] = 16'h0D50;
        ram[229] = 16'h2A8B;
        ram[230] = 16'h0470;
        ram[231] = 16'h2E2F;
        ram[232] = 16'h117B;
        ram[233] = 16'h0F65;
        ram[234] = 16'h15D4;
        ram[235] = 16'h1522;
        ram[236] = 16'h1747;
        ram[237] = 16'h270C;
        ram[238] = 16'h27C3;
        ram[239] = 16'h0D04;
        ram[240] = 16'h0D41;
        ram[241] = 16'h1457;
        ram[242] = 16'h046B;
        ram[243] = 16'h16C8;
        ram[244] = 16'h0179;
        ram[245] = 16'h0798;
        ram[246] = 16'h107E;
        ram[247] = 16'h0288;
        ram[248] = 16'h2580;
        ram[249] = 16'h00D8;
        ram[250] = 16'h0C80;
        ram[251] = 16'h0048;
        ram[252] = 16'h142B;
        ram[253] = 16'h0018;
        ram[254] = 16'h06B9;
        ram[255] = 16'h0008;
        ram[256] = 16'h123E;
        ram[257] = 16'h1003;
        ram[258] = 16'h1615;
        ram[259] = 16'h2557;
        ram[260] = 16'h275D;
        ram[261] = 16'h2C73;
        ram[262] = 16'h0D1F;
        ram[263] = 16'h0ED1;
        ram[264] = 16'h1460;
        ram[265] = 16'h24F1;
        ram[266] = 16'h16CB;
        ram[267] = 16'h2C51;
        ram[268] = 16'h0799;
        ram[269] = 16'h1EC6;
        ram[270] = 16'h2289;
        ram[271] = 16'h0A42;
        ram[272] = 16'h0B83;
        ram[273] = 16'h236C;
        ram[274] = 16'h23D7;
        ram[275] = 16'h1BCF;
        ram[276] = 16'h2BF3;
        ram[277] = 16'h0945;
        ram[278] = 16'h2EA7;
        ram[279] = 16'h0317;
        ram[280] = 16'h0F8D;
        ram[281] = 16'h1108;
        ram[282] = 16'h052F;
        ram[283] = 16'h25AE;
        ram[284] = 16'h21BB;
        ram[285] = 16'h2C90;
        ram[286] = 16'h2B3F;
        ram[287] = 16'h1EDB;
        ram[288] = 16'h2E6B;
        ram[289] = 16'h0A49;
        ram[290] = 16'h0F79;
        ram[291] = 16'h136E;
        ram[292] = 16'h2529;
        ram[293] = 16'h067A;
        ram[294] = 16'h0C63;
        ram[295] = 16'h1229;
        ram[296] = 16'h0421;
        ram[297] = 16'h160E;
        ram[298] = 16'h2161;
        ram[299] = 16'h075A;
        ram[300] = 16'h2B21;
        ram[301] = 16'h2274;
        ram[302] = 16'h2E61;
        ram[303] = 16'h0B7C;
        ram[304] = 16'h1F76;
        ram[305] = 16'h03D4;
        ram[306] = 16'h1A7D;
        ram[307] = 16'h1147;
        ram[308] = 16'h28D5;
        ram[309] = 16'h25C3;
        ram[310] = 16'h2D9D;
        ram[311] = 16'h2C97;
        ram[312] = 16'h2F35;
        ram[313] = 16'h0EDD;
        ram[314] = 16'h2FBD;
        ram[315] = 16'h24F5;
        ram[316] = 16'h1FEA;
        ram[317] = 16'h1C52;
        ram[318] = 16'h2AA4;
        ram[319] = 16'h1971;
        ram[320] = 16'h1E37;
        ram[321] = 16'h087B;
        ram[322] = 16'h2A13;
        ram[323] = 16'h12D4;
        ram[324] = 16'h2E07;
        ram[325] = 16'h1647;
        ram[326] = 16'h1F58;
        ram[327] = 16'h076D;
        ram[328] = 16'h1A73;
        ram[329] = 16'h127A;
        ram[330] = 16'h08D1;
        ram[331] = 16'h1629;
        ram[332] = 16'h22F1;
        ram[333] = 16'h0763;
        ram[334] = 16'h1BA6;
        ram[335] = 16'h2277;
        ram[336] = 16'h2938;
        ram[337] = 16'h0B7D;
        ram[338] = 16'h2DBE;
        ram[339] = 16'h23D5;
        ram[340] = 16'h2F40;
        ram[341] = 16'h1BF2;
        ram[342] = 16'h0FC0;
        ram[343] = 16'h1951;
        ram[344] = 16'h0540;
        ram[345] = 16'h2871;
        ram[346] = 16'h01C0;
        ram[347] = 16'h0D7B;
        ram[348] = 16'h2096;
        ram[349] = 16'h247F;
        ram[350] = 16'h1ADD;
        ram[351] = 16'h2C2B;
        ram[352] = 16'h28F5;
        ram[353] = 16'h0EB9;
        ram[354] = 16'h0DA7;
        ram[355] = 16'h24E9;
        ram[356] = 16'h048D;
        ram[357] = 16'h1C4E;
        ram[358] = 16'h2185;
        ram[359] = 16'h2970;
        ram[360] = 16'h2B2D;
        ram[361] = 16'h0DD0;
        ram[362] = 16'h2E65;
        ram[363] = 16'h149B;
        ram[364] = 16'h0F77;
        ram[365] = 16'h26DF;
        ram[366] = 16'h1528;
        ram[367] = 16'h0CF5;
        ram[368] = 16'h270E;
        ram[369] = 16'h1452;
        ram[370] = 16'h1D05;
        ram[371] = 16'h06C6;
        ram[372] = 16'h29AD;
        ram[373] = 16'h0242;
        ram[374] = 16'h2DE5;
        ram[375] = 16'h10C1;
        ram[376] = 16'h2F4D;
        ram[377] = 16'h1596;
        ram[378] = 16'h2FC5;
        ram[379] = 16'h0732;
        ram[380] = 16'h2FED;
        ram[381] = 16'h0266;
        ram[382] = 16'h1FFA;
        ram[383] = 16'h10CD;
        ram[384] = 16'h1AA9;
        ram[385] = 16'h159A;
        ram[386] = 16'h08E3;
        ram[387] = 16'h2734;
        ram[388] = 16'h22F7;
        ram[389] = 16'h2D12;
        ram[390] = 16'h1BA8;
        ram[391] = 16'h0F06;
        ram[392] = 16'h0938;
        ram[393] = 16'h0502;
        ram[394] = 16'h1313;
        ram[395] = 16'h21AC;
        ram[396] = 16'h165C;
        ram[397] = 16'h2B3A;
        ram[398] = 16'h0774;
        ram[399] = 16'h1E69;
        ram[400] = 16'h027C;
        ram[401] = 16'h0A23;
        ram[402] = 16'h00D4;
        ram[403] = 16'h0361;
        ram[404] = 16'h1047;
        ram[405] = 16'h2121;
        ram[406] = 16'h056D;
        ram[407] = 16'h0B0B;
        ram[408] = 16'h01CF;
        ram[409] = 16'h23AF;
        ram[410] = 16'h209B;
        ram[411] = 16'h0BE5;
        ram[412] = 16'h2ADF;
        ram[413] = 16'h03F7;
        ram[414] = 16'h2E4B;
        ram[415] = 16'h2153;
        ram[416] = 16'h2F6F;
        ram[417] = 16'h1B1C;
        ram[418] = 16'h1FD0;
        ram[419] = 16'h290A;
        ram[420] = 16'h1A9B;
        ram[421] = 16'h0DAE;
        ram[422] = 16'h28DF;
        ram[423] = 16'h2490;
        ram[424] = 16'h1DA0;
        ram[425] = 16'h0C30;
        ram[426] = 16'h09E0;
        ram[427] = 16'h0410;
        ram[428] = 16'h134B;
        ram[429] = 16'h115B;
        ram[430] = 16'h266F;
        ram[431] = 16'h05C9;
        ram[432] = 16'h1CD0;
        ram[433] = 16'h11EE;
        ram[434] = 16'h199B;
        ram[435] = 16'h05FA;
        ram[436] = 16'h0889;
        ram[437] = 16'h01FE;
        ram[438] = 16'h22D9;
        ram[439] = 16'h00AA;
        ram[440] = 16'h1B9E;
        ram[441] = 16'h1039;
        ram[442] = 16'h1935;
        ram[443] = 16'h2569;
        ram[444] = 16'h0867;
        ram[445] = 16'h2C79;
        ram[446] = 16'h02CD;
        ram[447] = 16'h0ED3;
        ram[448] = 16'h00EF;
        ram[449] = 16'h04F1;
        ram[450] = 16'h1050;
        ram[451] = 16'h11A6;
        ram[452] = 16'h0570;
        ram[453] = 16'h05E2;
        ram[454] = 16'h01D0;
        ram[455] = 16'h01F6;
        ram[456] = 16'h109B;
        ram[457] = 16'h20A8;
        ram[458] = 16'h0589;
        ram[459] = 16'h1AE3;
        ram[460] = 16'h21D9;
        ram[461] = 16'h28F7;
        ram[462] = 16'h2B49;
        ram[463] = 16'h1DA8;
        ram[464] = 16'h1E6E;
        ram[465] = 16'h19E3;
        ram[466] = 16'h1A25;
        ram[467] = 16'h08A1;
        ram[468] = 16'h08B7;
        ram[469] = 16'h22E1;
        ram[470] = 16'h12E8;
        ram[471] = 16'h2BA1;
        ram[472] = 16'h264E;
        ram[473] = 16'h0E8B;
        ram[474] = 16'h1CC5;
        ram[475] = 16'h04D9;
        ram[476] = 16'h0997;
        ram[477] = 16'h119E;
        ram[478] = 16'h2333;
        ram[479] = 16'h25E0;
        ram[480] = 16'h1BBC;
        ram[481] = 16'h0CA0;
        ram[482] = 16'h193F;
        ram[483] = 16'h2436;
        ram[484] = 16'h286B;
        ram[485] = 16'h0C12;
        ram[486] = 16'h0D79;
        ram[487] = 16'h0406;
        ram[488] = 16'h147E;
        ram[489] = 16'h2158;
        ram[490] = 16'h16D5;
        ram[491] = 16'h2B1E;
        ram[492] = 16'h279D;
        ram[493] = 16'h2E60;
        ram[494] = 16'h2D35;
        ram[495] = 16'h2F76;
        ram[496] = 16'h1F12;
        ram[497] = 16'h0FD2;
        ram[498] = 16'h2A5C;
        ram[499] = 16'h0546;
        ram[500] = 16'h1E1F;
        ram[501] = 16'h01C2;
        ram[502] = 16'h2A0B;
        ram[503] = 16'h0096;
        ram[504] = 16'h1E04;
        ram[505] = 16'h0032;
        ram[506] = 16'h2A02;
        ram[507] = 16'h1011;
        ram[508] = 16'h1E01;
        ram[509] = 16'h055B;
        ram[510] = 16'h2A01;
        ram[511] = 16'h01C9;
       end else begin
        ram[0] = 16'h0FEB;
        ram[1] = 16'h14C3;
        ram[2] = 16'h1F1D;
        ram[3] = 16'h1CCD;
        ram[4] = 16'h020A;
        ram[5] = 16'h2788;
        ram[6] = 16'h2343;
        ram[7] = 16'h13D7;
        ram[8] = 16'h0928;
        ram[9] = 16'h04FE;
        ram[10] = 16'h07B5;
        ram[11] = 16'h15C6;
        ram[12] = 16'h03FA;
        ram[13] = 16'h18DC;
        ram[14] = 16'h2BF0;
        ram[15] = 16'h2247;
        ram[16] = 16'h1D4C;
        ram[17] = 16'h1E8E;
        ram[18] = 16'h15A1;
        ram[19] = 16'h128D;
        ram[20] = 16'h2134;
        ram[21] = 16'h2F6E;
        ram[22] = 16'h1550;
        ram[23] = 16'h1EA0;
        ram[24] = 16'h1545;
        ram[25] = 16'h0F14;
        ram[26] = 16'h11B8;
        ram[27] = 16'h2BE7;
        ram[28] = 16'h181B;
        ram[29] = 16'h2117;
        ram[30] = 16'h0A7B;
        ram[31] = 16'h2B5B;
        ram[32] = 16'h2941;
        ram[33] = 16'h0190;
        ram[34] = 16'h17F9;
        ram[35] = 16'h1CAD;
        ram[36] = 16'h1527;
        ram[37] = 16'h21C6;
        ram[38] = 16'h17F8;
        ram[39] = 16'h16E6;
        ram[40] = 16'h1599;
        ram[41] = 16'h1456;
        ram[42] = 16'h0038;
        ram[43] = 16'h2382;
        ram[44] = 16'h2214;
        ram[45] = 16'h2D73;
        ram[46] = 16'h06A6;
        ram[47] = 16'h283E;
        ram[48] = 16'h14DB;
        ram[49] = 16'h1ABB;
        ram[50] = 16'h17CD;
        ram[51] = 16'h0E7E;
        ram[52] = 16'h013C;
        ram[53] = 16'h017E;
        ram[54] = 16'h2E2D;
        ram[55] = 16'h206D;
        ram[56] = 16'h2AB2;
        ram[57] = 16'h153B;
        ram[58] = 16'h2B1B;
        ram[59] = 16'h03CD;
        ram[60] = 16'h2063;
        ram[61] = 16'h2810;
        ram[62] = 16'h20DA;
        ram[63] = 16'h0782;
        ram[64] = 16'h2F41;
        ram[65] = 16'h2AD8;
        ram[66] = 16'h2800;
        ram[67] = 16'h1330;
        ram[68] = 16'h125A;
        ram[69] = 16'h13C1;
        ram[70] = 16'h1D55;
        ram[71] = 16'h228C;
        ram[72] = 16'h2267;
        ram[73] = 16'h2CEE;
        ram[74] = 16'h155C;
        ram[75] = 16'h03F2;
        ram[76] = 16'h23CA;
        ram[77] = 16'h1FB8;
        ram[78] = 16'h0B68;
        ram[79] = 16'h1479;
        ram[80] = 16'h17A7;
        ram[81] = 16'h22F9;
        ram[82] = 16'h02A5;
        ram[83] = 16'h16F2;
        ram[84] = 16'h0ACE;
        ram[85] = 16'h2AD6;
        ram[86] = 16'h2FCD;
        ram[87] = 16'h239B;
        ram[88] = 16'h2F6A;
        ram[89] = 16'h27B2;
        ram[90] = 16'h0F75;
        ram[91] = 16'h0B17;
        ram[92] = 16'h18EF;
        ram[93] = 16'h09C9;
        ram[94] = 16'h2E52;
        ram[95] = 16'h062B;
        ram[96] = 16'h2342;
        ram[97] = 16'h0E10;
        ram[98] = 16'h17BD;
        ram[99] = 16'h1210;
        ram[100] = 16'h2E5C;
        ram[101] = 16'h0FF0;
        ram[102] = 16'h17B4;
        ram[103] = 16'h0E12;
        ram[104] = 16'h025D;
        ram[105] = 16'h2703;
        ram[106] = 16'h01F8;
        ram[107] = 16'h1F8C;
        ram[108] = 16'h12AE;
        ram[109] = 16'h1903;
        ram[110] = 16'h0BD5;
        ram[111] = 16'h1A27;
        ram[112] = 16'h2BB0;
        ram[113] = 16'h008E;
        ram[114] = 16'h1631;
        ram[115] = 16'h226C;
        ram[116] = 16'h0B1C;
        ram[117] = 16'h0D6E;
        ram[118] = 16'h1F8D;
        ram[119] = 16'h03CF;
        ram[120] = 16'h003A;
        ram[121] = 16'h2F10;
        ram[122] = 16'h03EB;
        ram[123] = 16'h2235;
        ram[124] = 16'h0375;
        ram[125] = 16'h1889;
        ram[126] = 16'h07A4;
        ram[127] = 16'h1391;
        ram[128] = 16'h2FC1;
        ram[129] = 16'h0E48;
        ram[130] = 16'h2D56;
        ram[131] = 16'h2666;
        ram[132] = 16'h061E;
        ram[133] = 16'h1696;
        ram[134] = 16'h09C7;
        ram[135] = 16'h0B84;
        ram[136] = 16'h1B78;
        ram[137] = 16'h0EFA;
        ram[138] = 16'h171F;
        ram[139] = 16'h1151;
        ram[140] = 16'h0BEE;
        ram[141] = 16'h1A93;
        ram[142] = 16'h23CE;
        ram[143] = 16'h06D3;
        ram[144] = 16'h27E3;
        ram[145] = 16'h2BA9;
        ram[146] = 16'h10E2;
        ram[147] = 16'h07A6;
        ram[148] = 16'h039A;
        ram[149] = 16'h2E48;
        ram[150] = 16'h0FEF;
        ram[151] = 16'h2BDF;
        ram[152] = 16'h0FCE;
        ram[153] = 16'h2D3C;
        ram[154] = 16'h0527;
        ram[155] = 16'h23B3;
        ram[156] = 16'h1850;
        ram[157] = 16'h0343;
        ram[158] = 16'h1F71;
        ram[159] = 16'h220F;
        ram[160] = 16'h1BC1;
        ram[161] = 16'h04B0;
        ram[162] = 16'h17EA;
        ram[163] = 16'h2606;
        ram[164] = 16'h0F74;
        ram[165] = 16'h0550;
        ram[166] = 16'h17E7;
        ram[167] = 16'h14B1;
        ram[168] = 16'h10CA;
        ram[169] = 16'h0D01;
        ram[170] = 16'h00A8;
        ram[171] = 16'h0A84;
        ram[172] = 16'h063A;
        ram[173] = 16'h2857;
        ram[174] = 16'h13F2;
        ram[175] = 16'h18B8;
        ram[176] = 16'h0E90;
        ram[177] = 16'h2030;
        ram[178] = 16'h1766;
        ram[179] = 16'h2B7A;
        ram[180] = 16'h03B4;
        ram[181] = 16'h047A;
        ram[182] = 16'h2A85;
        ram[183] = 16'h0145;
        ram[184] = 16'h2014;
        ram[185] = 16'h0FB0;
        ram[186] = 16'h214F;
        ram[187] = 16'h0B67;
        ram[188] = 16'h0127;
        ram[189] = 16'h182E;
        ram[190] = 16'h028C;
        ram[191] = 16'h1686;
        ram[192] = 16'h2DC1;
        ram[193] = 16'h2086;
        ram[194] = 16'h17FE;
        ram[195] = 16'h098F;
        ram[196] = 16'h070D;
        ram[197] = 16'h0B42;
        ram[198] = 16'h27FE;
        ram[199] = 16'h07A2;
        ram[200] = 16'h0733;
        ram[201] = 16'h26C8;
        ram[202] = 16'h1013;
        ram[203] = 16'h0BD6;
        ram[204] = 16'h0B5C;
        ram[205] = 16'h2F27;
        ram[206] = 16'h2238;
        ram[207] = 16'h0D6A;
        ram[208] = 16'h16F4;
        ram[209] = 16'h08E9;
        ram[210] = 16'h07EF;
        ram[211] = 16'h14D5;
        ram[212] = 16'h206A;
        ram[213] = 16'h2080;
        ram[214] = 16'h2F65;
        ram[215] = 16'h0ACF;
        ram[216] = 16'h2E3C;
        ram[217] = 16'h1714;
        ram[218] = 16'h2E5F;
        ram[219] = 16'h2145;
        ram[220] = 16'h1ACC;
        ram[221] = 16'h1D5B;
        ram[222] = 16'h2AF4;
        ram[223] = 16'h1281;
        ram[224] = 16'h09C4;
        ram[225] = 16'h2A30;
        ram[226] = 16'h1736;
        ram[227] = 16'h062F;
        ram[228] = 16'h2B12;
        ram[229] = 16'h2FD0;
        ram[230] = 16'h171B;
        ram[231] = 16'h2A36;
        ram[232] = 16'h0717;
        ram[233] = 16'h1507;
        ram[234] = 16'h05E8;
        ram[235] = 16'h2EA3;
        ram[236] = 16'h0809;
        ram[237] = 16'h1B08;
        ram[238] = 16'h237F;
        ram[239] = 16'h1E74;
        ram[240] = 16'h230E;
        ram[241] = 16'h01AA;
        ram[242] = 16'h1292;
        ram[243] = 16'h0742;
        ram[244] = 16'h2154;
        ram[245] = 16'h284A;
        ram[246] = 16'h2EA6;
        ram[247] = 16'h0B6D;
        ram[248] = 16'h00AE;
        ram[249] = 16'h2D2E;
        ram[250] = 16'h0BC1;
        ram[251] = 16'h069D;
        ram[252] = 16'h0A5F;
        ram[253] = 16'h199A;
        ram[254] = 16'h16EC;
        ram[255] = 16'h0AB2;
        ram[256] = 16'h2E14;
        ram[257] = 16'h2001;
        ram[258] = 16'h26B4;
        ram[259] = 16'h1544;
        ram[260] = 16'h2A9F;
        ram[261] = 16'h0778;
        ram[262] = 16'h1F10;
        ram[263] = 16'h01B3;
        ram[264] = 16'h0194;
        ram[265] = 16'h1DDC;
        ram[266] = 16'h2BD8;
        ram[267] = 16'h27A2;
        ram[268] = 16'h1B64;
        ram[269] = 16'h2B71;
        ram[270] = 16'h2B4A;
        ram[271] = 16'h2351;
        ram[272] = 16'h25FB;
        ram[273] = 16'h088B;
        ram[274] = 16'h268B;
        ram[275] = 16'h186A;
        ram[276] = 16'h0E3E;
        ram[277] = 16'h267C;
        ram[278] = 16'h187B;
        ram[279] = 16'h0BAB;
        ram[280] = 16'h213D;
        ram[281] = 16'h036B;
        ram[282] = 16'h1370;
        ram[283] = 16'h29BA;
        ram[284] = 16'h1F45;
        ram[285] = 16'h13E0;
        ram[286] = 16'h1C6E;
        ram[287] = 16'h2C17;
        ram[288] = 16'h2407;
        ram[289] = 16'h001B;
        ram[290] = 16'h0EB3;
        ram[291] = 16'h2A61;
        ram[292] = 16'h2C08;
        ram[293] = 16'h1CEC;
        ram[294] = 16'h13DC;
        ram[295] = 16'h29A1;
        ram[296] = 16'h1FD2;
        ram[297] = 16'h126A;
        ram[298] = 16'h2F0F;
        ram[299] = 16'h2A00;
        ram[300] = 16'h0A76;
        ram[301] = 16'h0E78;
        ram[302] = 16'h0221;
        ram[303] = 16'h1C66;
        ram[304] = 16'h042B;
        ram[305] = 16'h13ED;
        ram[306] = 16'h01BA;
        ram[307] = 16'h0961;
        ram[308] = 16'h0186;
        ram[309] = 16'h2CFC;
        ram[310] = 16'h0EC2;
        ram[311] = 16'h2108;
        ram[312] = 16'h0415;
        ram[313] = 16'h24D6;
        ram[314] = 16'h2650;
        ram[315] = 16'h1394;
        ram[316] = 16'h24A1;
        ram[317] = 16'h19BF;
        ram[318] = 16'h2E9F;
        ram[319] = 16'h12FD;
        ram[320] = 16'h1EAC;
        ram[321] = 16'h0003;
        ram[322] = 16'h0C4D;
        ram[323] = 16'h2F61;
        ram[324] = 16'h2F90;
        ram[325] = 16'h1337;
        ram[326] = 16'h278B;
        ram[327] = 16'h0F4B;
        ram[328] = 16'h0E34;
        ram[329] = 16'h1CB7;
        ram[330] = 16'h0A90;
        ram[331] = 16'h14AB;
        ram[332] = 16'h067F;
        ram[333] = 16'h06F1;
        ram[334] = 16'h0592;
        ram[335] = 16'h1DD3;
        ram[336] = 16'h05CC;
        ram[337] = 16'h1CE2;
        ram[338] = 16'h0ADC;
        ram[339] = 16'h1BB6;
        ram[340] = 16'h202C;
        ram[341] = 16'h0A55;
        ram[342] = 16'h1C4F;
        ram[343] = 16'h0901;
        ram[344] = 16'h0B1F;
        ram[345] = 16'h1EC3;
        ram[346] = 16'h1EED;
        ram[347] = 16'h2783;
        ram[348] = 16'h2968;
        ram[349] = 16'h22DD;
        ram[350] = 16'h0FD9;
        ram[351] = 16'h0CC7;
        ram[352] = 16'h2439;
        ram[353] = 16'h00F3;
        ram[354] = 16'h2449;
        ram[355] = 16'h2D62;
        ram[356] = 16'h0C40;
        ram[357] = 16'h1447;
        ram[358] = 16'h22B9;
        ram[359] = 16'h26A2;
        ram[360] = 16'h2E5D;
        ram[361] = 16'h15B7;
        ram[362] = 16'h277F;
        ram[363] = 16'h29F9;
        ram[364] = 16'h2E25;
        ram[365] = 16'h2236;
        ram[366] = 16'h1329;
        ram[367] = 16'h0F91;
        ram[368] = 16'h2583;
        ram[369] = 16'h2352;
        ram[370] = 16'h0F8A;
        ram[371] = 16'h2468;
        ram[372] = 16'h0DB6;
        ram[373] = 16'h14D4;
        ram[374] = 16'h24D0;
        ram[375] = 16'h0942;
        ram[376] = 16'h24BD;
        ram[377] = 16'h2B80;
        ram[378] = 16'h08C9;
        ram[379] = 16'h2031;
        ram[380] = 16'h29A3;
        ram[381] = 16'h27B3;
        ram[382] = 16'h238F;
        ram[383] = 16'h1AE2;
        ram[384] = 16'h2A3A;
        ram[385] = 16'h0001;
        ram[386] = 16'h141A;
        ram[387] = 16'h0FCB;
        ram[388] = 16'h1FDB;
        ram[389] = 16'h1668;
        ram[390] = 16'h2D2F;
        ram[391] = 16'h0519;
        ram[392] = 16'h04BC;
        ram[393] = 16'h2993;
        ram[394] = 16'h2386;
        ram[395] = 16'h16E4;
        ram[396] = 16'h222B;
        ram[397] = 16'h2251;
        ram[398] = 16'h21DC;
        ram[399] = 16'h09F1;
        ram[400] = 16'h11EF;
        ram[401] = 16'h19A1;
        ram[402] = 16'h139F;
        ram[403] = 16'h193D;
        ram[404] = 16'h2ABA;
        ram[405] = 16'h1372;
        ram[406] = 16'h1970;
        ram[407] = 16'h2301;
        ram[408] = 16'h03B5;
        ram[409] = 16'h0A41;
        ram[410] = 16'h0A4F;
        ram[411] = 16'h1D2C;
        ram[412] = 16'h2DCE;
        ram[413] = 16'h0B9F;
        ram[414] = 16'h2549;
        ram[415] = 16'h2443;
        ram[416] = 16'h0C13;
        ram[417] = 16'h0051;
        ram[418] = 16'h2C19;
        ram[419] = 16'h1F21;
        ram[420] = 16'h2416;
        ram[421] = 16'h26C3;
        ram[422] = 16'h0B93;
        ram[423] = 16'h1CE1;
        ram[424] = 16'h2F75;
        ram[425] = 16'h073D;
        ram[426] = 16'h2D2B;
        ram[427] = 16'h1DFE;
        ram[428] = 16'h1F62;
        ram[429] = 16'h2B68;
        ram[430] = 16'h0663;
        ram[431] = 16'h2531;
        ram[432] = 16'h0C81;
        ram[433] = 16'h0BC6;
        ram[434] = 16'h052E;
        ram[435] = 16'h1C23;
        ram[436] = 16'h0492;
        ram[437] = 16'h26F2;
        ram[438] = 16'h2C46;
        ram[439] = 16'h0316;
        ram[440] = 16'h0C3F;
        ram[441] = 16'h0E80;
        ram[442] = 16'h12EE;
        ram[443] = 16'h0ABB;
        ram[444] = 16'h0DE1;
        ram[445] = 16'h1D3C;
        ram[446] = 16'h2BDB;
        ram[447] = 16'h08F6;
        ram[448] = 16'h2C03;
        ram[449] = 16'h0009;
        ram[450] = 16'h24E7;
        ram[451] = 16'h2E21;
        ram[452] = 16'h2EAE;
        ram[453] = 16'h09A4;
        ram[454] = 16'h169F;
        ram[455] = 16'h2DE1;
        ram[456] = 16'h2A9C;
        ram[457] = 16'h2624;
        ram[458] = 16'h1FB0;
        ram[459] = 16'h0E00;
        ram[460] = 16'h137D;
        ram[461] = 16'h14D3;
        ram[462] = 16'h10B6;
        ram[463] = 16'h2978;
        ram[464] = 16'h1164;
        ram[465] = 16'h26A5;
        ram[466] = 16'h2094;
        ram[467] = 16'h2321;
        ram[468] = 16'h0082;
        ram[469] = 16'h1EFF;
        ram[470] = 16'h24EC;
        ram[471] = 16'h1B03;
        ram[472] = 16'h215D;
        ram[473] = 16'h2C48;
        ram[474] = 16'h2CC6;
        ram[475] = 16'h1687;
        ram[476] = 16'h1C36;
        ram[477] = 16'h0895;
        ram[478] = 16'h2F8B;
        ram[479] = 16'h2655;
        ram[480] = 16'h0CA9;
        ram[481] = 16'h02D9;
        ram[482] = 16'h0CD9;
        ram[483] = 16'h2824;
        ram[484] = 16'h24C0;
        ram[485] = 16'h0CD4;
        ram[486] = 16'h0829;
        ram[487] = 16'h13E4;
        ram[488] = 16'h2B15;
        ram[489] = 16'h1124;
        ram[490] = 16'h167B;
        ram[491] = 16'h1DE9;
        ram[492] = 16'h2A6D;
        ram[493] = 16'h06A0;
        ram[494] = 16'h097A;
        ram[495] = 16'h2EB3;
        ram[496] = 16'h1087;
        ram[497] = 16'h09F4;
        ram[498] = 16'h2E9E;
        ram[499] = 16'h0D36;
        ram[500] = 16'h2922;
        ram[501] = 16'h0E7B;
        ram[502] = 16'h0E6E;
        ram[503] = 16'h1BC6;
        ram[504] = 16'h0E35;
        ram[505] = 16'h227E;
        ram[506] = 16'h1A5B;
        ram[507] = 16'h0091;
        ram[508] = 16'h1CE7;
        ram[509] = 16'h1717;
        ram[510] = 16'h0AAB;
        ram[511] = 16'h20A5;
       end
       */
    
    
endmodule