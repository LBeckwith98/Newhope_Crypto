`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07/13/2020 09:45:35 PM
// Design Name: 
// Module Name: bitrev_map
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module bitrev_mapfull(
    input [8:0] in_addr,
    output reg [8:0] out_addr
    );
    
    always @(*) begin
    case(in_addr)
        0: out_addr = 9'd0;
        1: out_addr = 9'd256;
        2: out_addr = 9'd128;
        3: out_addr = 9'd384;
        4: out_addr = 9'd64;
        5: out_addr = 9'd320;
        6: out_addr = 9'd192;
        7: out_addr = 9'd448;
        8: out_addr = 9'd32;
        9: out_addr = 9'd288;
        10: out_addr = 9'd160;
        11: out_addr = 9'd416;
        12: out_addr = 9'd96;
        13: out_addr = 9'd352;
        14: out_addr = 9'd224;
        15: out_addr = 9'd480;
        16: out_addr = 9'd16;
        17: out_addr = 9'd272;
        18: out_addr = 9'd144;
        19: out_addr = 9'd400;
        20: out_addr = 9'd80;
        21: out_addr = 9'd336;
        22: out_addr = 9'd208;
        23: out_addr = 9'd464;
        24: out_addr = 9'd48;
        25: out_addr = 9'd304;
        26: out_addr = 9'd176;
        27: out_addr = 9'd432;
        28: out_addr = 9'd112;
        29: out_addr = 9'd368;
        30: out_addr = 9'd240;
        31: out_addr = 9'd496;
        32: out_addr = 9'd8;
        33: out_addr = 9'd264;
        34: out_addr = 9'd136;
        35: out_addr = 9'd392;
        36: out_addr = 9'd72;
        37: out_addr = 9'd328;
        38: out_addr = 9'd200;
        39: out_addr = 9'd456;
        40: out_addr = 9'd40;
        41: out_addr = 9'd296;
        42: out_addr = 9'd168;
        43: out_addr = 9'd424;
        44: out_addr = 9'd104;
        45: out_addr = 9'd360;
        46: out_addr = 9'd232;
        47: out_addr = 9'd488;
        48: out_addr = 9'd24;
        49: out_addr = 9'd280;
        50: out_addr = 9'd152;
        51: out_addr = 9'd408;
        52: out_addr = 9'd88;
        53: out_addr = 9'd344;
        54: out_addr = 9'd216;
        55: out_addr = 9'd472;
        56: out_addr = 9'd56;
        57: out_addr = 9'd312;
        58: out_addr = 9'd184;
        59: out_addr = 9'd440;
        60: out_addr = 9'd120;
        61: out_addr = 9'd376;
        62: out_addr = 9'd248;
        63: out_addr = 9'd504;
        64: out_addr = 9'd4;
        65: out_addr = 9'd260;
        66: out_addr = 9'd132;
        67: out_addr = 9'd388;
        68: out_addr = 9'd68;
        69: out_addr = 9'd324;
        70: out_addr = 9'd196;
        71: out_addr = 9'd452;
        72: out_addr = 9'd36;
        73: out_addr = 9'd292;
        74: out_addr = 9'd164;
        75: out_addr = 9'd420;
        76: out_addr = 9'd100;
        77: out_addr = 9'd356;
        78: out_addr = 9'd228;
        79: out_addr = 9'd484;
        80: out_addr = 9'd20;
        81: out_addr = 9'd276;
        82: out_addr = 9'd148;
        83: out_addr = 9'd404;
        84: out_addr = 9'd84;
        85: out_addr = 9'd340;
        86: out_addr = 9'd212;
        87: out_addr = 9'd468;
        88: out_addr = 9'd52;
        89: out_addr = 9'd308;
        90: out_addr = 9'd180;
        91: out_addr = 9'd436;
        92: out_addr = 9'd116;
        93: out_addr = 9'd372;
        94: out_addr = 9'd244;
        95: out_addr = 9'd500;
        96: out_addr = 9'd12;
        97: out_addr = 9'd268;
        98: out_addr = 9'd140;
        99: out_addr = 9'd396;
        100: out_addr = 9'd76;
        101: out_addr = 9'd332;
        102: out_addr = 9'd204;
        103: out_addr = 9'd460;
        104: out_addr = 9'd44;
        105: out_addr = 9'd300;
        106: out_addr = 9'd172;
        107: out_addr = 9'd428;
        108: out_addr = 9'd108;
        109: out_addr = 9'd364;
        110: out_addr = 9'd236;
        111: out_addr = 9'd492;
        112: out_addr = 9'd28;
        113: out_addr = 9'd284;
        114: out_addr = 9'd156;
        115: out_addr = 9'd412;
        116: out_addr = 9'd92;
        117: out_addr = 9'd348;
        118: out_addr = 9'd220;
        119: out_addr = 9'd476;
        120: out_addr = 9'd60;
        121: out_addr = 9'd316;
        122: out_addr = 9'd188;
        123: out_addr = 9'd444;
        124: out_addr = 9'd124;
        125: out_addr = 9'd380;
        126: out_addr = 9'd252;
        127: out_addr = 9'd508;
        128: out_addr = 9'd2;
        129: out_addr = 9'd258;
        130: out_addr = 9'd130;
        131: out_addr = 9'd386;
        132: out_addr = 9'd66;
        133: out_addr = 9'd322;
        134: out_addr = 9'd194;
        135: out_addr = 9'd450;
        136: out_addr = 9'd34;
        137: out_addr = 9'd290;
        138: out_addr = 9'd162;
        139: out_addr = 9'd418;
        140: out_addr = 9'd98;
        141: out_addr = 9'd354;
        142: out_addr = 9'd226;
        143: out_addr = 9'd482;
        144: out_addr = 9'd18;
        145: out_addr = 9'd274;
        146: out_addr = 9'd146;
        147: out_addr = 9'd402;
        148: out_addr = 9'd82;
        149: out_addr = 9'd338;
        150: out_addr = 9'd210;
        151: out_addr = 9'd466;
        152: out_addr = 9'd50;
        153: out_addr = 9'd306;
        154: out_addr = 9'd178;
        155: out_addr = 9'd434;
        156: out_addr = 9'd114;
        157: out_addr = 9'd370;
        158: out_addr = 9'd242;
        159: out_addr = 9'd498;
        160: out_addr = 9'd10;
        161: out_addr = 9'd266;
        162: out_addr = 9'd138;
        163: out_addr = 9'd394;
        164: out_addr = 9'd74;
        165: out_addr = 9'd330;
        166: out_addr = 9'd202;
        167: out_addr = 9'd458;
        168: out_addr = 9'd42;
        169: out_addr = 9'd298;
        170: out_addr = 9'd170;
        171: out_addr = 9'd426;
        172: out_addr = 9'd106;
        173: out_addr = 9'd362;
        174: out_addr = 9'd234;
        175: out_addr = 9'd490;
        176: out_addr = 9'd26;
        177: out_addr = 9'd282;
        178: out_addr = 9'd154;
        179: out_addr = 9'd410;
        180: out_addr = 9'd90;
        181: out_addr = 9'd346;
        182: out_addr = 9'd218;
        183: out_addr = 9'd474;
        184: out_addr = 9'd58;
        185: out_addr = 9'd314;
        186: out_addr = 9'd186;
        187: out_addr = 9'd442;
        188: out_addr = 9'd122;
        189: out_addr = 9'd378;
        190: out_addr = 9'd250;
        191: out_addr = 9'd506;
        192: out_addr = 9'd6;
        193: out_addr = 9'd262;
        194: out_addr = 9'd134;
        195: out_addr = 9'd390;
        196: out_addr = 9'd70;
        197: out_addr = 9'd326;
        198: out_addr = 9'd198;
        199: out_addr = 9'd454;
        200: out_addr = 9'd38;
        201: out_addr = 9'd294;
        202: out_addr = 9'd166;
        203: out_addr = 9'd422;
        204: out_addr = 9'd102;
        205: out_addr = 9'd358;
        206: out_addr = 9'd230;
        207: out_addr = 9'd486;
        208: out_addr = 9'd22;
        209: out_addr = 9'd278;
        210: out_addr = 9'd150;
        211: out_addr = 9'd406;
        212: out_addr = 9'd86;
        213: out_addr = 9'd342;
        214: out_addr = 9'd214;
        215: out_addr = 9'd470;
        216: out_addr = 9'd54;
        217: out_addr = 9'd310;
        218: out_addr = 9'd182;
        219: out_addr = 9'd438;
        220: out_addr = 9'd118;
        221: out_addr = 9'd374;
        222: out_addr = 9'd246;
        223: out_addr = 9'd502;
        224: out_addr = 9'd14;
        225: out_addr = 9'd270;
        226: out_addr = 9'd142;
        227: out_addr = 9'd398;
        228: out_addr = 9'd78;
        229: out_addr = 9'd334;
        230: out_addr = 9'd206;
        231: out_addr = 9'd462;
        232: out_addr = 9'd46;
        233: out_addr = 9'd302;
        234: out_addr = 9'd174;
        235: out_addr = 9'd430;
        236: out_addr = 9'd110;
        237: out_addr = 9'd366;
        238: out_addr = 9'd238;
        239: out_addr = 9'd494;
        240: out_addr = 9'd30;
        241: out_addr = 9'd286;
        242: out_addr = 9'd158;
        243: out_addr = 9'd414;
        244: out_addr = 9'd94;
        245: out_addr = 9'd350;
        246: out_addr = 9'd222;
        247: out_addr = 9'd478;
        248: out_addr = 9'd62;
        249: out_addr = 9'd318;
        250: out_addr = 9'd190;
        251: out_addr = 9'd446;
        252: out_addr = 9'd126;
        253: out_addr = 9'd382;
        254: out_addr = 9'd254;
        255: out_addr = 9'd510;
        256: out_addr = 9'd1;
        257: out_addr = 9'd257;
        258: out_addr = 9'd129;
        259: out_addr = 9'd385;
        260: out_addr = 9'd65;
        261: out_addr = 9'd321;
        262: out_addr = 9'd193;
        263: out_addr = 9'd449;
        264: out_addr = 9'd33;
        265: out_addr = 9'd289;
        266: out_addr = 9'd161;
        267: out_addr = 9'd417;
        268: out_addr = 9'd97;
        269: out_addr = 9'd353;
        270: out_addr = 9'd225;
        271: out_addr = 9'd481;
        272: out_addr = 9'd17;
        273: out_addr = 9'd273;
        274: out_addr = 9'd145;
        275: out_addr = 9'd401;
        276: out_addr = 9'd81;
        277: out_addr = 9'd337;
        278: out_addr = 9'd209;
        279: out_addr = 9'd465;
        280: out_addr = 9'd49;
        281: out_addr = 9'd305;
        282: out_addr = 9'd177;
        283: out_addr = 9'd433;
        284: out_addr = 9'd113;
        285: out_addr = 9'd369;
        286: out_addr = 9'd241;
        287: out_addr = 9'd497;
        288: out_addr = 9'd9;
        289: out_addr = 9'd265;
        290: out_addr = 9'd137;
        291: out_addr = 9'd393;
        292: out_addr = 9'd73;
        293: out_addr = 9'd329;
        294: out_addr = 9'd201;
        295: out_addr = 9'd457;
        296: out_addr = 9'd41;
        297: out_addr = 9'd297;
        298: out_addr = 9'd169;
        299: out_addr = 9'd425;
        300: out_addr = 9'd105;
        301: out_addr = 9'd361;
        302: out_addr = 9'd233;
        303: out_addr = 9'd489;
        304: out_addr = 9'd25;
        305: out_addr = 9'd281;
        306: out_addr = 9'd153;
        307: out_addr = 9'd409;
        308: out_addr = 9'd89;
        309: out_addr = 9'd345;
        310: out_addr = 9'd217;
        311: out_addr = 9'd473;
        312: out_addr = 9'd57;
        313: out_addr = 9'd313;
        314: out_addr = 9'd185;
        315: out_addr = 9'd441;
        316: out_addr = 9'd121;
        317: out_addr = 9'd377;
        318: out_addr = 9'd249;
        319: out_addr = 9'd505;
        320: out_addr = 9'd5;
        321: out_addr = 9'd261;
        322: out_addr = 9'd133;
        323: out_addr = 9'd389;
        324: out_addr = 9'd69;
        325: out_addr = 9'd325;
        326: out_addr = 9'd197;
        327: out_addr = 9'd453;
        328: out_addr = 9'd37;
        329: out_addr = 9'd293;
        330: out_addr = 9'd165;
        331: out_addr = 9'd421;
        332: out_addr = 9'd101;
        333: out_addr = 9'd357;
        334: out_addr = 9'd229;
        335: out_addr = 9'd485;
        336: out_addr = 9'd21;
        337: out_addr = 9'd277;
        338: out_addr = 9'd149;
        339: out_addr = 9'd405;
        340: out_addr = 9'd85;
        341: out_addr = 9'd341;
        342: out_addr = 9'd213;
        343: out_addr = 9'd469;
        344: out_addr = 9'd53;
        345: out_addr = 9'd309;
        346: out_addr = 9'd181;
        347: out_addr = 9'd437;
        348: out_addr = 9'd117;
        349: out_addr = 9'd373;
        350: out_addr = 9'd245;
        351: out_addr = 9'd501;
        352: out_addr = 9'd13;
        353: out_addr = 9'd269;
        354: out_addr = 9'd141;
        355: out_addr = 9'd397;
        356: out_addr = 9'd77;
        357: out_addr = 9'd333;
        358: out_addr = 9'd205;
        359: out_addr = 9'd461;
        360: out_addr = 9'd45;
        361: out_addr = 9'd301;
        362: out_addr = 9'd173;
        363: out_addr = 9'd429;
        364: out_addr = 9'd109;
        365: out_addr = 9'd365;
        366: out_addr = 9'd237;
        367: out_addr = 9'd493;
        368: out_addr = 9'd29;
        369: out_addr = 9'd285;
        370: out_addr = 9'd157;
        371: out_addr = 9'd413;
        372: out_addr = 9'd93;
        373: out_addr = 9'd349;
        374: out_addr = 9'd221;
        375: out_addr = 9'd477;
        376: out_addr = 9'd61;
        377: out_addr = 9'd317;
        378: out_addr = 9'd189;
        379: out_addr = 9'd445;
        380: out_addr = 9'd125;
        381: out_addr = 9'd381;
        382: out_addr = 9'd253;
        383: out_addr = 9'd509;
        384: out_addr = 9'd3;
        385: out_addr = 9'd259;
        386: out_addr = 9'd131;
        387: out_addr = 9'd387;
        388: out_addr = 9'd67;
        389: out_addr = 9'd323;
        390: out_addr = 9'd195;
        391: out_addr = 9'd451;
        392: out_addr = 9'd35;
        393: out_addr = 9'd291;
        394: out_addr = 9'd163;
        395: out_addr = 9'd419;
        396: out_addr = 9'd99;
        397: out_addr = 9'd355;
        398: out_addr = 9'd227;
        399: out_addr = 9'd483;
        400: out_addr = 9'd19;
        401: out_addr = 9'd275;
        402: out_addr = 9'd147;
        403: out_addr = 9'd403;
        404: out_addr = 9'd83;
        405: out_addr = 9'd339;
        406: out_addr = 9'd211;
        407: out_addr = 9'd467;
        408: out_addr = 9'd51;
        409: out_addr = 9'd307;
        410: out_addr = 9'd179;
        411: out_addr = 9'd435;
        412: out_addr = 9'd115;
        413: out_addr = 9'd371;
        414: out_addr = 9'd243;
        415: out_addr = 9'd499;
        416: out_addr = 9'd11;
        417: out_addr = 9'd267;
        418: out_addr = 9'd139;
        419: out_addr = 9'd395;
        420: out_addr = 9'd75;
        421: out_addr = 9'd331;
        422: out_addr = 9'd203;
        423: out_addr = 9'd459;
        424: out_addr = 9'd43;
        425: out_addr = 9'd299;
        426: out_addr = 9'd171;
        427: out_addr = 9'd427;
        428: out_addr = 9'd107;
        429: out_addr = 9'd363;
        430: out_addr = 9'd235;
        431: out_addr = 9'd491;
        432: out_addr = 9'd27;
        433: out_addr = 9'd283;
        434: out_addr = 9'd155;
        435: out_addr = 9'd411;
        436: out_addr = 9'd91;
        437: out_addr = 9'd347;
        438: out_addr = 9'd219;
        439: out_addr = 9'd475;
        440: out_addr = 9'd59;
        441: out_addr = 9'd315;
        442: out_addr = 9'd187;
        443: out_addr = 9'd443;
        444: out_addr = 9'd123;
        445: out_addr = 9'd379;
        446: out_addr = 9'd251;
        447: out_addr = 9'd507;
        448: out_addr = 9'd7;
        449: out_addr = 9'd263;
        450: out_addr = 9'd135;
        451: out_addr = 9'd391;
        452: out_addr = 9'd71;
        453: out_addr = 9'd327;
        454: out_addr = 9'd199;
        455: out_addr = 9'd455;
        456: out_addr = 9'd39;
        457: out_addr = 9'd295;
        458: out_addr = 9'd167;
        459: out_addr = 9'd423;
        460: out_addr = 9'd103;
        461: out_addr = 9'd359;
        462: out_addr = 9'd231;
        463: out_addr = 9'd487;
        464: out_addr = 9'd23;
        465: out_addr = 9'd279;
        466: out_addr = 9'd151;
        467: out_addr = 9'd407;
        468: out_addr = 9'd87;
        469: out_addr = 9'd343;
        470: out_addr = 9'd215;
        471: out_addr = 9'd471;
        472: out_addr = 9'd55;
        473: out_addr = 9'd311;
        474: out_addr = 9'd183;
        475: out_addr = 9'd439;
        476: out_addr = 9'd119;
        477: out_addr = 9'd375;
        478: out_addr = 9'd247;
        479: out_addr = 9'd503;
        480: out_addr = 9'd15;
        481: out_addr = 9'd271;
        482: out_addr = 9'd143;
        483: out_addr = 9'd399;
        484: out_addr = 9'd79;
        485: out_addr = 9'd335;
        486: out_addr = 9'd207;
        487: out_addr = 9'd463;
        488: out_addr = 9'd47;
        489: out_addr = 9'd303;
        490: out_addr = 9'd175;
        491: out_addr = 9'd431;
        492: out_addr = 9'd111;
        493: out_addr = 9'd367;
        494: out_addr = 9'd239;
        495: out_addr = 9'd495;
        496: out_addr = 9'd31;
        497: out_addr = 9'd287;
        498: out_addr = 9'd159;
        499: out_addr = 9'd415;
        500: out_addr = 9'd95;
        501: out_addr = 9'd351;
        502: out_addr = 9'd223;
        503: out_addr = 9'd479;
        504: out_addr = 9'd63;
        505: out_addr = 9'd319;
        506: out_addr = 9'd191;
        507: out_addr = 9'd447;
        508: out_addr = 9'd127;
        509: out_addr = 9'd383;
        510: out_addr = 9'd255;
        511: out_addr = 9'd511;
    endcase
    end
endmodule